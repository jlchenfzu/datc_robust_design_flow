VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x2_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.136 0.144 0.944 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.828 0.108 1.224 0.18 ;
        RECT 0.828 0.736 0.9 0.972 ;
        RECT 0.828 0.108 0.9 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.72 0.972 ;
      RECT 0.648 0.108 0.72 0.972 ;
      RECT 0.648 0.504 0.812 0.576 ;
      RECT 0.28 0.108 0.352 0.344 ;
      RECT 0.28 0.108 0.72 0.18 ;
  END
END AND2x2_ASAP7_75t_R

MACRO AND2x4_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x4_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.112 1.008 0.6 ;
        RECT 0.288 0.112 1.008 0.184 ;
        RECT 0.288 0.112 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.428 0.576 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.24 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.924 0.972 ;
      RECT 0.72 0.256 0.792 0.972 ;
      RECT 0.716 0.728 1.224 0.8 ;
      RECT 1.152 0.484 1.224 0.8 ;
      RECT 0.46 0.256 0.792 0.328 ;
  END
END AND2x4_ASAP7_75t_R

MACRO AND2x6_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x6_ASAP7_75t_R 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.112 1.008 0.6 ;
        RECT 0.288 0.112 1.008 0.184 ;
        RECT 0.288 0.112 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.428 0.576 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 2.216 0.972 ;
        RECT 1.24 0.108 2.216 0.18 ;
        RECT 1.8 0.108 1.872 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.924 0.972 ;
      RECT 0.72 0.256 0.792 0.972 ;
      RECT 0.716 0.728 1.224 0.8 ;
      RECT 1.152 0.484 1.224 0.8 ;
      RECT 0.46 0.256 0.792 0.328 ;
  END
END AND2x6_ASAP7_75t_R

MACRO AND3x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x1_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.732 1.224 0.804 ;
        RECT 1.152 0.304 1.224 0.804 ;
        RECT 1.044 0.304 1.224 0.376 ;
        RECT 1.044 0.732 1.116 0.94 ;
        RECT 1.044 0.136 1.116 0.376 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.936 0.972 ;
      RECT 0.864 0.108 0.936 0.972 ;
      RECT 0.864 0.504 1.052 0.576 ;
      RECT 0.16 0.108 0.936 0.18 ;
  END
END AND3x1_ASAP7_75t_R

MACRO AND3x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x2_ASAP7_75t_R 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.044 0.108 1.44 0.18 ;
        RECT 1.044 0.736 1.116 0.972 ;
        RECT 1.044 0.108 1.116 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.936 0.972 ;
      RECT 0.864 0.108 0.936 0.972 ;
      RECT 0.864 0.504 1.136 0.576 ;
      RECT 0.16 0.108 0.936 0.18 ;
  END
END AND3x2_ASAP7_75t_R

MACRO AND3x4_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x4_ASAP7_75t_R 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.756 2.596 0.828 ;
        RECT 2.448 0.396 2.596 0.468 ;
        RECT 2.448 0.396 2.52 0.828 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.756 2.164 0.828 ;
        RECT 2.016 0.396 2.164 0.468 ;
        RECT 2.016 0.396 2.088 0.828 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.92 0.972 ;
        RECT 0.072 0.108 0.92 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.04 0.9 2.984 0.972 ;
      RECT 2.912 0.108 2.984 0.972 ;
      RECT 1.04 0.168 1.112 0.972 ;
      RECT 0.872 0.504 1.112 0.576 ;
      RECT 2.536 0.108 2.984 0.18 ;
      RECT 1.888 0.252 2.804 0.324 ;
      RECT 1.24 0.108 2.216 0.18 ;
  END
END AND3x4_ASAP7_75t_R

MACRO AND4x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x1_ASAP7_75t_R 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.136 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.136 0.792 0.8 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.136 1.008 0.656 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.196 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.24 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 1.008 0.972 ;
      RECT 0.936 0.756 1.008 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.936 0.756 1.224 0.828 ;
      RECT 1.152 0.48 1.224 0.828 ;
      RECT 0.072 0.108 0.34 0.18 ;
  END
END AND4x1_ASAP7_75t_R

MACRO AND4x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x2_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.136 1.224 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.136 1.008 0.8 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.136 0.792 0.656 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.488 0.972 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.9 1.656 0.972 ;
      RECT 1.584 0.108 1.656 0.972 ;
      RECT 0.612 0.756 0.684 0.972 ;
      RECT 0.396 0.756 0.684 0.828 ;
      RECT 0.396 0.476 0.468 0.828 ;
      RECT 1.456 0.108 1.656 0.18 ;
  END
END AND4x2_ASAP7_75t_R

MACRO AOI211x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211x1_ASAP7_75t_R 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.504 0.916 0.576 ;
        RECT 0.72 0.756 0.892 0.828 ;
        RECT 0.72 0.252 0.88 0.324 ;
        RECT 0.72 0.252 0.792 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.492 0.576 ;
        RECT 0.072 0.136 0.144 0.944 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.612 1.768 0.684 ;
        RECT 1.584 0.252 1.768 0.324 ;
        RECT 1.584 0.252 1.656 0.684 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.504 2.216 0.576 ;
        RECT 2.016 0.252 2.2 0.324 ;
        RECT 2.016 0.252 2.088 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.076 0.756 2.52 0.828 ;
        RECT 2.448 0.108 2.52 0.828 ;
        RECT 0.364 0.108 2.52 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.9 1.224 0.972 ;
      RECT 1.152 0.756 1.224 0.972 ;
      RECT 1.152 0.756 1.796 0.828 ;
      RECT 1.444 0.9 2.432 0.972 ;
  END
END AOI211x1_ASAP7_75t_R

MACRO AOI211xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.36 0.576 ;
        RECT 0.072 0.28 0.144 0.8 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.16 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.704 0.972 ;
  END
END AOI211xp5_ASAP7_75t_R

MACRO AOI21x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21x1_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.252 1.224 0.656 ;
        RECT 0.504 0.252 1.224 0.324 ;
        RECT 0.504 0.252 0.576 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.76 0.5 1.024 0.572 ;
        RECT 0.76 0.396 0.908 0.684 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.756 1.44 0.828 ;
        RECT 1.368 0.464 1.44 0.828 ;
        RECT 0.288 0.28 0.36 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.476 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.072 0.108 1.656 0.18 ;
        RECT 0.072 0.9 0.252 0.972 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.9 1.332 0.972 ;
  END
END AOI21x1_ASAP7_75t_R

MACRO AOI21xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21xp33_ASAP7_75t_R 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.5 0.38 0.572 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.428 0.108 1.008 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.684 0.972 ;
  END
END AOI21xp33_ASAP7_75t_R

MACRO AOI21xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.5 0.38 0.572 ;
        RECT 0.072 0.136 0.144 0.8 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.568 0.108 1.008 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.684 0.972 ;
  END
END AOI21xp5_ASAP7_75t_R

MACRO AOI221x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221x1_ASAP7_75t_R 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.612 0.868 0.684 ;
        RECT 0.72 0.108 0.792 0.684 ;
        RECT 0.644 0.108 0.792 0.18 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.504 0.596 0.576 ;
        RECT 0.212 0.612 0.36 0.684 ;
        RECT 0.288 0.108 0.36 0.684 ;
        RECT 0.212 0.108 0.36 0.18 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.324 1.3 0.396 ;
        RECT 1.076 0.612 1.224 0.684 ;
        RECT 1.152 0.324 1.224 0.684 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.612 1.948 0.684 ;
        RECT 1.8 0.324 1.872 0.684 ;
        RECT 1.564 0.504 1.872 0.576 ;
        RECT 1.724 0.324 1.872 0.396 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.504 2.544 0.576 ;
        RECT 2.156 0.756 2.304 0.828 ;
        RECT 2.232 0.324 2.304 0.828 ;
        RECT 2.156 0.324 2.304 0.396 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.536 0.756 2.952 0.828 ;
        RECT 2.88 0.18 2.952 0.828 ;
        RECT 1.024 0.18 2.952 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.24 0.9 2.864 0.972 ;
      RECT 0.16 0.756 2 0.828 ;
  END
END AOI221x1_ASAP7_75t_R

MACRO AOI221xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.136 1.224 0.656 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.92 0.18 ;
        RECT 0.072 0.756 0.492 0.828 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.804 0.756 1.356 0.828 ;
      RECT 0.16 0.9 0.704 0.972 ;
  END
END AOI221xp5_ASAP7_75t_R

MACRO AOI222xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222xp33_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.136 1.872 0.8 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 1.596 0.18 ;
        RECT 0.072 0.756 0.488 0.828 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.368 0.9 1.872 0.972 ;
      RECT 1.368 0.756 1.44 0.972 ;
      RECT 0.808 0.756 1.44 0.828 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END AOI222xp33_ASAP7_75t_R

MACRO AOI22x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22x1_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.612 1.516 0.684 ;
        RECT 1.368 0.396 1.516 0.468 ;
        RECT 1.368 0.396 1.44 0.684 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.724 0.612 1.872 0.684 ;
        RECT 1.8 0.252 1.872 0.684 ;
        RECT 1.152 0.252 1.872 0.324 ;
        RECT 1.152 0.252 1.224 0.608 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.756 0.792 0.828 ;
        RECT 0.72 0.396 0.792 0.828 ;
        RECT 0.644 0.396 0.792 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.616 ;
        RECT 0.288 0.252 1.008 0.324 ;
        RECT 0.288 0.756 0.436 0.828 ;
        RECT 0.288 0.252 0.36 0.828 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.236 0.756 2.088 0.828 ;
        RECT 2.016 0.108 2.088 0.828 ;
        RECT 0.152 0.108 2.088 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 2 0.972 ;
  END
END AOI22x1_ASAP7_75t_R

MACRO AOI22xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22xp33_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.136 0.36 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.592 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END AOI22xp33_ASAP7_75t_R

MACRO AOI22xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.28 0.576 0.828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.592 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END AOI22xp5_ASAP7_75t_R

MACRO BUFx10_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx10_ASAP7_75t_R 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.9 2.952 0.972 ;
        RECT 2.88 0.108 2.952 0.972 ;
        RECT 0.796 0.108 2.952 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 2.756 0.576 ;
      RECT 0.364 0.108 0.576 0.18 ;
  END
END BUFx10_ASAP7_75t_R

MACRO BUFx12_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx12_ASAP7_75t_R 0 0 ;
  SIZE 3.456 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.456 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.9 3.384 0.972 ;
        RECT 3.312 0.108 3.384 0.972 ;
        RECT 0.796 0.108 3.384 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 3.2 0.576 ;
      RECT 0.376 0.108 0.576 0.18 ;
  END
END BUFx12_ASAP7_75t_R

MACRO BUFx12f_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx12f_ASAP7_75t_R 0 0 ;
  SIZE 3.888 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.136 0.144 0.944 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.888 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.888 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 3.816 0.972 ;
        RECT 3.744 0.108 3.816 0.972 ;
        RECT 1.24 0.108 3.816 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 1.116 0.972 ;
      RECT 1.044 0.108 1.116 0.972 ;
      RECT 1.044 0.504 1.244 0.576 ;
      RECT 0.376 0.108 1.116 0.18 ;
  END
END BUFx12f_ASAP7_75t_R

MACRO BUFx16f_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx16f_ASAP7_75t_R 0 0 ;
  SIZE 4.752 BY 1.08 ;
  SYMMETRY X Y ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.752 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.752 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 4.68 0.972 ;
        RECT 4.608 0.108 4.68 0.972 ;
        RECT 1.24 0.108 4.68 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.936 0.504 4.496 0.576 ;
      RECT 0.376 0.108 1.008 0.18 ;
      RECT 0.072 0.136 0.144 0.944 ;
  END
END BUFx16f_ASAP7_75t_R

MACRO BUFx24_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx24_ASAP7_75t_R 0 0 ;
  SIZE 6.48 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 6.48 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.48 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 6.408 0.972 ;
        RECT 6.336 0.108 6.408 0.972 ;
        RECT 1.24 0.108 6.408 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.936 0.504 6.212 0.576 ;
      RECT 0.376 0.108 1.008 0.18 ;
  END
END BUFx24_ASAP7_75t_R

MACRO BUFx2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx2_ASAP7_75t_R 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.58 0.108 1.008 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 0.812 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUFx2_ASAP7_75t_R

MACRO BUFx3_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx3_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.58 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 1.04 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUFx3_ASAP7_75t_R

MACRO BUFx4_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4_ASAP7_75t_R 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 1.428 0.972 ;
        RECT 1.356 0.108 1.428 0.972 ;
        RECT 0.58 0.108 1.428 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 1.256 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUFx4_ASAP7_75t_R

MACRO BUFx4f_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4f_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.392 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.796 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 1.468 0.576 ;
      RECT 0.364 0.108 0.576 0.18 ;
  END
END BUFx4f_ASAP7_75t_R

MACRO BUFx5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx5_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.58 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 1.472 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUFx5_ASAP7_75t_R

MACRO BUFx6f_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx6f_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.136 0.144 0.944 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 2.088 0.972 ;
        RECT 2.016 0.108 2.088 0.972 ;
        RECT 0.808 0.108 2.088 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 1.892 0.576 ;
      RECT 0.376 0.108 0.576 0.18 ;
  END
END BUFx6f_ASAP7_75t_R

MACRO BUFx8_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx8_ASAP7_75t_R 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.392 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 2.52 0.972 ;
        RECT 2.448 0.108 2.52 0.972 ;
        RECT 0.808 0.108 2.52 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 2.324 0.576 ;
      RECT 0.364 0.108 0.576 0.18 ;
  END
END BUFx8_ASAP7_75t_R

MACRO DFFHQx4_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQx4_ASAP7_75t_R 0 0 ;
  SIZE 5.4 BY 1.08 ;
  SYMMETRY X Y ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.656 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.424 ;
        RECT 0.396 0.136 0.468 0.424 ;
        RECT 0.288 0.656 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.504 1.16 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5 0.9 5.332 0.972 ;
        RECT 5.252 0.108 5.332 0.972 ;
        RECT 4.5 0.108 5.332 0.18 ;
        RECT 4.5 0.804 4.572 0.972 ;
        RECT 4.5 0.108 4.572 0.276 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.4 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.4 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.048 0.9 4.392 0.972 ;
      RECT 4.32 0.108 4.392 0.972 ;
      RECT 4.32 0.508 4.7 0.58 ;
      RECT 4.048 0.108 4.392 0.18 ;
      RECT 3.4 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.096 0.108 3.168 0.476 ;
      RECT 3.096 0.108 3.816 0.18 ;
      RECT 2.752 0.896 2.952 0.968 ;
      RECT 2.88 0.108 2.952 0.968 ;
      RECT 2.88 0.612 3.6 0.684 ;
      RECT 3.528 0.468 3.6 0.684 ;
      RECT 3.312 0.468 3.384 0.684 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 2.304 0.9 2.52 0.972 ;
      RECT 2.448 0.324 2.52 0.972 ;
      RECT 1.984 0.324 2.52 0.396 ;
      RECT 2.34 0.18 2.412 0.396 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.324 0.56 ;
      RECT 1.672 0.108 1.872 0.18 ;
      RECT 1.26 0.504 1.332 0.812 ;
      RECT 1.26 0.504 1.468 0.576 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.576 0.188 0.648 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.96 0.488 4.032 0.668 ;
      RECT 2.664 0.404 2.736 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.668 ;
      RECT 0.568 0.424 0.64 0.668 ;
    LAYER M2 ;
      RECT 3.508 0.576 4.052 0.648 ;
      RECT 0.076 0.576 2.756 0.648 ;
      RECT 0.7 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 3.96 0.576 4.032 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.664 0.576 2.736 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.26 0.72 1.332 0.792 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.568 0.576 0.64 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END DFFHQx4_ASAP7_75t_R

MACRO INVx11_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx11_ASAP7_75t_R 0 0 ;
  SIZE 2.808 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.808 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 2.736 0.972 ;
        RECT 2.664 0.108 2.736 0.972 ;
        RECT 0.376 0.108 2.736 0.18 ;
    END
  END Y
END INVx11_ASAP7_75t_R

MACRO INVx13_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx13_ASAP7_75t_R 0 0 ;
  SIZE 3.24 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.24 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 3.168 0.972 ;
        RECT 3.096 0.108 3.168 0.972 ;
        RECT 0.376 0.108 3.168 0.18 ;
    END
  END Y
END INVx13_ASAP7_75t_R

MACRO INVx1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx1_ASAP7_75t_R 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.576 0.972 ;
        RECT 0.504 0.108 0.576 0.972 ;
        RECT 0.376 0.108 0.576 0.18 ;
    END
  END Y
END INVx1_ASAP7_75t_R

MACRO INVx2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx2_ASAP7_75t_R 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.376 0.108 0.792 0.18 ;
    END
  END Y
END INVx2_ASAP7_75t_R

MACRO INVx3_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx3_ASAP7_75t_R 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.376 0.108 1.008 0.18 ;
    END
  END Y
END INVx3_ASAP7_75t_R

MACRO INVx4_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx4_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.376 0.108 1.224 0.18 ;
    END
  END Y
END INVx4_ASAP7_75t_R

MACRO INVx5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx5_ASAP7_75t_R 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 0.376 0.108 1.44 0.18 ;
    END
  END Y
END INVx5_ASAP7_75t_R

MACRO INVx6_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx6_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.376 0.108 1.656 0.18 ;
    END
  END Y
END INVx6_ASAP7_75t_R

MACRO INVx8_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx8_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 2.088 0.972 ;
        RECT 2.016 0.108 2.088 0.972 ;
        RECT 0.376 0.108 2.088 0.18 ;
    END
  END Y
END INVx8_ASAP7_75t_R

MACRO INVxp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVxp33_ASAP7_75t_R 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.136 0.144 0.944 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.576 0.972 ;
        RECT 0.504 0.108 0.576 0.972 ;
        RECT 0.376 0.108 0.576 0.18 ;
    END
  END Y
END INVxp33_ASAP7_75t_R

MACRO INVxp67_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVxp67_ASAP7_75t_R 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.136 0.144 0.944 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.576 0.972 ;
        RECT 0.504 0.108 0.576 0.972 ;
        RECT 0.376 0.108 0.576 0.18 ;
    END
  END Y
END INVxp67_ASAP7_75t_R

MACRO NAND2x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.26 0.144 0.944 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.224 0.972 ;
        RECT 1.152 0.252 1.224 0.972 ;
        RECT 0.808 0.252 1.224 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END NAND2x1_ASAP7_75t_R

MACRO NAND2x1p5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1p5_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.136 0.144 0.944 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 1.028 0.576 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 1.044 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.252 1.352 0.324 ;
      RECT 0.376 0.108 0.9 0.18 ;
  END
END NAND2x1p5_ASAP7_75t_R

MACRO NAND2x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x2_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.968 0.756 1.116 0.828 ;
        RECT 1.044 0.424 1.116 0.828 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.396 1.872 0.708 ;
        RECT 1.288 0.396 1.872 0.468 ;
        RECT 1.288 0.252 1.36 0.468 ;
        RECT 0.8 0.252 1.36 0.324 ;
        RECT 0.288 0.396 0.872 0.468 ;
        RECT 0.8 0.252 0.872 0.468 ;
        RECT 0.288 0.756 0.436 0.828 ;
        RECT 0.288 0.396 0.36 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 2.088 0.972 ;
        RECT 2.016 0.252 2.088 0.972 ;
        RECT 1.672 0.252 2.088 0.324 ;
        RECT 0.072 0.252 0.488 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 2 0.18 ;
  END
END NAND2x2_ASAP7_75t_R

MACRO NAND2xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp33_ASAP7_75t_R 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.572 0.108 0.792 0.18 ;
    END
  END Y
END NAND2xp33_ASAP7_75t_R

MACRO NAND2xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp5_ASAP7_75t_R 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.424 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.572 0.108 0.792 0.18 ;
    END
  END Y
END NAND2xp5_ASAP7_75t_R

MACRO NAND2xp67_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp67_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.5 0.38 0.572 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 0.756 1.008 0.828 ;
        RECT 0.936 0.424 1.008 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.9 1.224 0.972 ;
        RECT 1.152 0.252 1.224 0.972 ;
        RECT 0.808 0.252 1.224 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END NAND2xp67_ASAP7_75t_R

MACRO NAND3x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x1_ASAP7_75t_R 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.608 0.72 1.872 0.792 ;
        RECT 1.8 0.432 1.872 0.792 ;
        RECT 1.6 0.432 1.872 0.504 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.972 0.72 1.224 0.792 ;
        RECT 1.152 0.432 1.224 0.792 ;
        RECT 0.984 0.432 1.224 0.504 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.244 0.412 0.316 0.812 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 2.304 0.972 ;
        RECT 2.232 0.252 2.304 0.972 ;
        RECT 1.672 0.252 2.304 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.024 0.108 2 0.18 ;
      RECT 0.376 0.252 1.352 0.324 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END NAND3x1_ASAP7_75t_R

MACRO NAND3x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x2_ASAP7_75t_R 0 0 ;
  SIZE 4.32 BY 1.08 ;
  SYMMETRY X Y ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.352 0.756 2.972 0.828 ;
        RECT 2.9 0.424 2.972 0.828 ;
        RECT 1.352 0.424 1.424 0.828 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.188 0.424 2.26 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.32 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 4.248 0.972 ;
        RECT 4.176 0.252 4.248 0.972 ;
        RECT 3.616 0.252 4.248 0.324 ;
        RECT 0.072 0.252 0.704 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.676 0.72 3.632 0.792 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 3.464 0.756 3.612 0.828 ;
      RECT 3.54 0.432 3.612 0.828 ;
      RECT 0.696 0.756 0.844 0.828 ;
      RECT 0.696 0.424 0.768 0.828 ;
      RECT 2.968 0.108 3.944 0.18 ;
      RECT 1.024 0.252 3.296 0.324 ;
      RECT 1.672 0.108 2.648 0.18 ;
      RECT 0.376 0.108 1.352 0.18 ;
    LAYER V1 ;
      RECT 3.54 0.72 3.612 0.792 ;
      RECT 0.696 0.72 0.768 0.792 ;
  END
END NAND3x2_ASAP7_75t_R

MACRO NAND3xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3xp33_ASAP7_75t_R 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.136 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.136 0.792 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.704 0.972 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
END NAND3xp33_ASAP7_75t_R

MACRO NAND4xp25_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4xp25_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.136 0.792 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.136 0.576 0.8 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.136 0.36 0.8 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.16 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 1.024 0.108 1.224 0.18 ;
    END
  END Y
END NAND4xp25_ASAP7_75t_R

MACRO NAND4xp75_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4xp75_ASAP7_75t_R 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.424 2.52 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.404 2.196 0.476 ;
        RECT 2.124 0.28 2.196 0.476 ;
        RECT 2.016 0.404 2.088 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.404 1.224 0.8 ;
        RECT 0.828 0.404 1.224 0.476 ;
        RECT 0.828 0.28 0.9 0.476 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.228 0.972 ;
        RECT 0.072 0.108 0.228 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 2.952 0.972 ;
        RECT 2.88 0.252 2.952 0.972 ;
        RECT 2.32 0.252 2.952 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.648 0.108 2.664 0.18 ;
      RECT 1.024 0.252 1.996 0.324 ;
      RECT 0.368 0.108 1.36 0.18 ;
  END
END NAND4xp75_ASAP7_75t_R

MACRO NOR2x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 0.92 0.576 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.376 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END NOR2x1_ASAP7_75t_R

MACRO NOR2x1p5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1p5_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 1.028 0.576 ;
        RECT 0.504 0.252 0.652 0.324 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.376 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.756 1.352 0.828 ;
      RECT 0.376 0.9 0.9 0.972 ;
  END
END NOR2x1p5_ASAP7_75t_R

MACRO NOR2x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x2_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.252 1.116 0.656 ;
        RECT 0.968 0.252 1.116 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.288 0.612 1.872 0.684 ;
        RECT 1.8 0.372 1.872 0.684 ;
        RECT 0.8 0.756 1.36 0.828 ;
        RECT 1.288 0.612 1.36 0.828 ;
        RECT 0.8 0.612 0.872 0.828 ;
        RECT 0.288 0.612 0.872 0.684 ;
        RECT 0.288 0.252 0.436 0.324 ;
        RECT 0.288 0.252 0.36 0.684 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.756 2.088 0.828 ;
        RECT 2.016 0.108 2.088 0.828 ;
        RECT 0.072 0.108 2.088 0.18 ;
        RECT 0.072 0.756 0.488 0.828 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 2 0.972 ;
  END
END NOR2x2_ASAP7_75t_R

MACRO NOR2xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2xp33_ASAP7_75t_R 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.572 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.376 0.108 0.792 0.18 ;
    END
  END Y
END NOR2xp33_ASAP7_75t_R

MACRO NOR2xp67_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2xp67_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.508 0.38 0.58 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 1.028 0.576 ;
        RECT 0.504 0.252 0.652 0.324 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.592 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END NOR2xp67_ASAP7_75t_R

MACRO NOR3x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x1_ASAP7_75t_R 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.612 1.872 0.684 ;
        RECT 1.8 0.252 1.872 0.684 ;
        RECT 1.584 0.252 1.872 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.612 1.224 0.684 ;
        RECT 1.152 0.252 1.224 0.684 ;
        RECT 0.936 0.252 1.224 0.324 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.36 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.756 2.304 0.828 ;
        RECT 2.232 0.108 2.304 0.828 ;
        RECT 0.808 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.024 0.9 2 0.972 ;
      RECT 0.376 0.756 1.352 0.828 ;
      RECT 0.16 0.9 0.704 0.972 ;
  END
END NOR3x1_ASAP7_75t_R

MACRO NOR3x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x2_ASAP7_75t_R 0 0 ;
  SIZE 4.32 BY 1.08 ;
  SYMMETRY X Y ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9 0.252 2.972 0.656 ;
        RECT 1.352 0.252 2.972 0.324 ;
        RECT 1.352 0.252 1.424 0.656 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.188 0.424 2.26 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.32 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.616 0.756 4.248 0.828 ;
        RECT 4.176 0.108 4.248 0.828 ;
        RECT 0.072 0.108 4.248 0.18 ;
        RECT 0.072 0.756 0.704 0.828 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.676 0.288 3.632 0.36 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 3.54 0.252 3.612 0.648 ;
      RECT 3.464 0.252 3.612 0.324 ;
      RECT 0.696 0.252 0.768 0.656 ;
      RECT 0.696 0.252 0.844 0.324 ;
      RECT 2.968 0.9 3.944 0.972 ;
      RECT 1.024 0.756 3.296 0.828 ;
      RECT 1.672 0.9 2.648 0.972 ;
      RECT 0.376 0.9 1.352 0.972 ;
    LAYER V1 ;
      RECT 3.54 0.288 3.612 0.36 ;
      RECT 0.696 0.288 0.768 0.36 ;
  END
END NOR3x2_ASAP7_75t_R

MACRO NOR3xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3xp33_ASAP7_75t_R 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.944 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.944 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.704 0.18 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
END NOR3xp33_ASAP7_75t_R

MACRO NOR4xp25_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4xp25_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.944 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.944 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.944 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.16 0.108 1.224 0.18 ;
    END
  END Y
END NOR4xp25_ASAP7_75t_R

MACRO NOR4xp75_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4xp75_ASAP7_75t_R 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.28 2.52 0.656 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.124 0.604 2.196 0.8 ;
        RECT 2.016 0.604 2.196 0.676 ;
        RECT 2.016 0.28 2.088 0.676 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.604 1.224 0.676 ;
        RECT 1.152 0.28 1.224 0.676 ;
        RECT 0.828 0.604 0.9 0.8 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.228 0.972 ;
        RECT 0.072 0.108 0.228 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.32 0.756 2.952 0.828 ;
        RECT 2.88 0.108 2.952 0.828 ;
        RECT 0.376 0.108 2.952 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.648 0.9 2.664 0.972 ;
      RECT 1.024 0.756 1.996 0.828 ;
      RECT 0.368 0.9 1.36 0.972 ;
  END
END NOR4xp75_ASAP7_75t_R

MACRO OAI211xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.36 0.576 ;
        RECT 0.072 0.28 0.144 0.8 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.16 0.9 1.224 0.972 ;
        RECT 1.152 0.252 1.224 0.972 ;
        RECT 0.396 0.252 1.224 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END OAI211xp5_ASAP7_75t_R

MACRO OAI21x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21x1_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.756 1.224 0.828 ;
        RECT 1.152 0.424 1.224 0.828 ;
        RECT 0.504 0.424 0.576 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.76 0.508 1.024 0.58 ;
        RECT 0.76 0.396 0.908 0.684 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.252 1.44 0.616 ;
        RECT 0.288 0.252 1.44 0.324 ;
        RECT 0.288 0.252 0.36 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 1.476 0.108 1.656 0.18 ;
        RECT 0.072 0.108 0.252 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.108 1.332 0.18 ;
  END
END OAI21x1_ASAP7_75t_R

MACRO OAI21xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21xp33_ASAP7_75t_R 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.28 0.144 0.944 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.812 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.9 1.008 0.972 ;
        RECT 0.936 0.252 1.008 0.972 ;
        RECT 0.396 0.252 1.008 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END OAI21xp33_ASAP7_75t_R

MACRO OAI21xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.28 0.144 0.944 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.812 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.684 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.9 1.008 0.972 ;
        RECT 0.936 0.252 1.008 0.972 ;
        RECT 0.396 0.252 1.008 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END OAI21xp5_ASAP7_75t_R

MACRO OAI221xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.944 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.424 0.36 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.92 0.972 ;
        RECT 0.072 0.252 0.492 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.804 0.252 1.356 0.324 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END OAI221xp5_ASAP7_75t_R

MACRO OAI222xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222xp33_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.424 0.36 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.8 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.8 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 2.088 0.972 ;
        RECT 2.016 0.22 2.088 0.972 ;
        RECT 0.072 0.252 0.488 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.252 1.44 0.324 ;
      RECT 1.368 0.108 1.44 0.324 ;
      RECT 1.368 0.108 1.872 0.18 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END OAI222xp33_ASAP7_75t_R

MACRO OAI22x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22x1_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.612 1.516 0.684 ;
        RECT 1.368 0.396 1.516 0.468 ;
        RECT 1.368 0.396 1.44 0.684 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.756 1.872 0.828 ;
        RECT 1.8 0.396 1.872 0.828 ;
        RECT 1.724 0.396 1.872 0.468 ;
        RECT 1.152 0.472 1.224 0.828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.612 0.792 0.684 ;
        RECT 0.72 0.252 0.792 0.684 ;
        RECT 0.644 0.252 0.792 0.324 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.756 1.008 0.828 ;
        RECT 0.936 0.464 1.008 0.828 ;
        RECT 0.288 0.252 0.436 0.324 ;
        RECT 0.288 0.252 0.36 0.828 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.152 0.9 2.088 0.972 ;
        RECT 2.016 0.252 2.088 0.972 ;
        RECT 1.236 0.252 2.088 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 2 0.18 ;
  END
END OAI22x1_ASAP7_75t_R

MACRO OAI22xp33_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22xp33_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.424 0.36 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.9 1.1 0.972 ;
        RECT 0.936 0.28 1.008 0.972 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.704 0.972 ;
        RECT 0.072 0.252 0.468 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END OAI22xp33_ASAP7_75t_R

MACRO OAI22xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.424 0.36 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.9 1.1 0.972 ;
        RECT 0.936 0.28 1.008 0.972 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.656 ;
        RECT 0.604 0.252 0.792 0.324 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.704 0.972 ;
        RECT 0.072 0.252 0.468 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END OAI22xp5_ASAP7_75t_R

MACRO OR2x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x2_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.828 0.108 1.224 0.18 ;
        RECT 0.828 0.736 0.9 0.972 ;
        RECT 0.828 0.108 0.9 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.744 0.972 ;
      RECT 0.672 0.108 0.744 0.972 ;
      RECT 0.672 0.504 0.908 0.576 ;
      RECT 0.376 0.108 0.744 0.18 ;
  END
END OR2x2_ASAP7_75t_R

MACRO OR2x4_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x4_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.828 0.108 1.656 0.18 ;
        RECT 1.26 0.736 1.332 0.972 ;
        RECT 1.26 0.108 1.332 0.344 ;
        RECT 0.828 0.736 0.9 0.972 ;
        RECT 0.828 0.108 0.9 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.748 0.972 ;
      RECT 0.676 0.108 0.748 0.972 ;
      RECT 0.676 0.504 0.908 0.576 ;
      RECT 0.376 0.108 0.748 0.18 ;
  END
END OR2x4_ASAP7_75t_R

MACRO OR2x6_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x6_ASAP7_75t_R 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.252 0.576 0.488 ;
        RECT 0.072 0.252 0.576 0.324 ;
        RECT 0.072 0.252 0.144 0.944 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.612 1.008 0.684 ;
        RECT 0.936 0.484 1.008 0.684 ;
        RECT 0.288 0.424 0.36 0.944 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.9 2.52 0.972 ;
        RECT 2.448 0.108 2.52 0.972 ;
        RECT 1.24 0.108 2.52 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.592 0.756 1.224 0.828 ;
      RECT 1.152 0.28 1.224 0.828 ;
      RECT 0.936 0.28 1.224 0.352 ;
      RECT 0.936 0.108 1.008 0.352 ;
      RECT 0.376 0.108 1.008 0.18 ;
  END
END OR2x6_ASAP7_75t_R

MACRO OR3x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x1_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.732 1.224 0.804 ;
        RECT 1.152 0.304 1.224 0.804 ;
        RECT 1.044 0.304 1.224 0.376 ;
        RECT 1.044 0.732 1.116 0.94 ;
        RECT 1.044 0.136 1.116 0.376 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.936 0.972 ;
      RECT 0.864 0.108 0.936 0.972 ;
      RECT 0.864 0.504 1.048 0.576 ;
      RECT 0.16 0.108 0.936 0.18 ;
  END
END OR3x1_ASAP7_75t_R

MACRO OR3x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x2_ASAP7_75t_R 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.044 0.108 1.44 0.18 ;
        RECT 1.044 0.736 1.116 0.972 ;
        RECT 1.044 0.108 1.116 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.96 0.972 ;
      RECT 0.888 0.108 0.96 0.972 ;
      RECT 0.888 0.504 1.136 0.576 ;
      RECT 0.16 0.108 0.96 0.18 ;
  END
END OR3x2_ASAP7_75t_R

MACRO OR3x4_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x4_ASAP7_75t_R 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.044 0.108 1.872 0.18 ;
        RECT 1.476 0.736 1.548 0.972 ;
        RECT 1.476 0.108 1.548 0.344 ;
        RECT 1.044 0.736 1.116 0.972 ;
        RECT 1.044 0.108 1.116 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.964 0.972 ;
      RECT 0.892 0.108 0.964 0.972 ;
      RECT 0.892 0.504 1.136 0.576 ;
      RECT 0.16 0.108 0.964 0.18 ;
  END
END OR3x4_ASAP7_75t_R

MACRO OR4x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4x1_ASAP7_75t_R 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.944 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.944 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.944 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.24 0.9 1.44 0.972 ;
      RECT 1.368 0.108 1.44 0.972 ;
      RECT 0.288 0.264 0.36 0.608 ;
      RECT 0.288 0.264 0.468 0.336 ;
      RECT 0.396 0.108 0.468 0.336 ;
      RECT 0.396 0.108 1.44 0.18 ;
  END
END OR4x1_ASAP7_75t_R

MACRO OR4x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4x2_ASAP7_75t_R 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.944 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.944 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.944 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.488 0.972 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.456 0.9 1.656 0.972 ;
      RECT 1.584 0.108 1.656 0.972 ;
      RECT 0.396 0.252 0.468 0.596 ;
      RECT 0.396 0.252 0.684 0.324 ;
      RECT 0.612 0.108 0.684 0.324 ;
      RECT 0.612 0.108 1.656 0.18 ;
  END
END OR4x2_ASAP7_75t_R

MACRO TIEHIx1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHIx1_ASAP7_75t_R 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  PIN H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.972 ;
    END
  END H
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.072 0.512 0.38 0.584 ;
      RECT 0.072 0.108 0.144 0.584 ;
      RECT 0.072 0.108 0.272 0.18 ;
      RECT 0.268 0.28 0.376 0.352 ;
  END
END TIEHIx1_ASAP7_75t_R

MACRO TIELOx1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELOx1_ASAP7_75t_R 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  PIN L
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.268 0.728 0.576 0.8 ;
        RECT 0.504 0.108 0.576 0.8 ;
        RECT 0.376 0.108 0.576 0.18 ;
    END
  END L
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 0.272 0.972 ;
      RECT 0.072 0.496 0.144 0.972 ;
      RECT 0.072 0.496 0.38 0.568 ;
  END
END TIELOx1_ASAP7_75t_R

MACRO XNOR2x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x1_ASAP7_75t_R 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.22 0.504 1.46 0.576 ;
        RECT 1.22 0.268 1.292 0.576 ;
        RECT 0.852 0.268 1.292 0.34 ;
        RECT 0.852 0.108 0.924 0.34 ;
        RECT 0.072 0.108 0.924 0.18 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.108 0.144 0.944 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.9 2.448 0.972 ;
        RECT 1.8 0.308 1.872 0.972 ;
        RECT 1.672 0.308 1.872 0.38 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.484 0.72 2.324 0.792 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 2.104 0.756 2.304 0.828 ;
      RECT 2.232 0.484 2.304 0.828 ;
      RECT 0.368 0.9 0.772 0.972 ;
      RECT 0.696 0.756 0.772 0.972 ;
      RECT 0.696 0.756 1.656 0.828 ;
      RECT 1.584 0.484 1.656 0.828 ;
      RECT 0.696 0.328 0.768 0.972 ;
      RECT 0.428 0.756 0.576 0.828 ;
      RECT 0.504 0.484 0.576 0.828 ;
      RECT 1.024 0.108 2.432 0.18 ;
      RECT 2.016 0.28 2.088 0.608 ;
    LAYER M2 ;
      RECT 1.192 0.288 2.108 0.36 ;
    LAYER V1 ;
      RECT 2.232 0.72 2.304 0.792 ;
      RECT 2.016 0.288 2.088 0.36 ;
      RECT 1.22 0.288 1.292 0.36 ;
      RECT 0.504 0.72 0.576 0.792 ;
  END
END XNOR2x1_ASAP7_75t_R

MACRO XNOR2x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x2_ASAP7_75t_R 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.76 0.972 ;
        RECT 1.688 0.504 1.76 0.972 ;
        RECT 1.564 0.504 1.76 0.576 ;
        RECT 1.044 0.732 1.116 0.972 ;
        RECT 0.504 0.732 1.116 0.804 ;
        RECT 0.504 0.48 0.576 0.804 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.756 1.52 0.828 ;
        RECT 1.368 0.428 1.44 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.888 0.9 2.304 0.972 ;
        RECT 2.232 0.108 2.304 0.972 ;
        RECT 1.888 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 0.252 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 1.908 0.252 1.98 0.604 ;
      RECT 1.692 0.252 1.98 0.324 ;
      RECT 1.692 0.108 1.764 0.324 ;
      RECT 0.072 0.108 1.764 0.18 ;
      RECT 1.208 0.252 1.28 0.78 ;
      RECT 0.288 0.252 0.36 0.596 ;
      RECT 0.288 0.252 1.568 0.324 ;
      RECT 0.396 0.9 0.92 0.972 ;
  END
END XNOR2x2_ASAP7_75t_R

MACRO XNOR2xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.252 1.44 0.656 ;
        RECT 0.828 0.252 1.44 0.324 ;
        RECT 0.828 0.108 0.9 0.324 ;
        RECT 0.288 0.108 0.9 0.18 ;
        RECT 0.288 0.108 0.36 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.692 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.72 0.972 ;
      RECT 0.648 0.3 0.72 0.972 ;
      RECT 0.648 0.756 1.656 0.828 ;
      RECT 1.584 0.484 1.656 0.828 ;
      RECT 1.044 0.108 1.548 0.18 ;
  END
END XNOR2xp5_ASAP7_75t_R

MACRO XOR2x1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x1_ASAP7_75t_R 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.22 0.504 1.46 0.576 ;
        RECT 0.852 0.74 1.292 0.812 ;
        RECT 1.22 0.504 1.292 0.812 ;
        RECT 0.072 0.9 0.924 0.972 ;
        RECT 0.852 0.74 0.924 0.972 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.136 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.108 2.448 0.18 ;
        RECT 1.672 0.7 1.872 0.772 ;
        RECT 1.8 0.108 1.872 0.772 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.484 0.288 2.324 0.36 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 2.232 0.252 2.304 0.596 ;
      RECT 2.104 0.252 2.304 0.324 ;
      RECT 0.696 0.108 0.768 0.752 ;
      RECT 1.584 0.252 1.656 0.596 ;
      RECT 0.696 0.252 1.656 0.324 ;
      RECT 0.696 0.108 0.772 0.324 ;
      RECT 0.368 0.108 0.772 0.18 ;
      RECT 0.504 0.252 0.576 0.596 ;
      RECT 0.428 0.252 0.576 0.324 ;
      RECT 1.024 0.9 2.432 0.972 ;
      RECT 2.016 0.472 2.088 0.8 ;
    LAYER M2 ;
      RECT 1.192 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 2.232 0.288 2.304 0.36 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.22 0.72 1.292 0.792 ;
      RECT 0.504 0.288 0.576 0.36 ;
  END
END XOR2x1_ASAP7_75t_R

MACRO XOR2x2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x2_ASAP7_75t_R 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.252 1.52 0.324 ;
        RECT 1.368 0.252 1.44 0.652 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.688 0.108 1.76 0.652 ;
        RECT 1.564 0.504 1.76 0.576 ;
        RECT 1.044 0.108 1.76 0.18 ;
        RECT 0.504 0.276 1.116 0.348 ;
        RECT 1.044 0.108 1.116 0.348 ;
        RECT 0.504 0.276 0.576 0.6 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.888 0.9 2.304 0.972 ;
        RECT 2.232 0.108 2.304 0.972 ;
        RECT 1.888 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 1.764 0.972 ;
      RECT 1.692 0.756 1.764 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 1.692 0.756 1.98 0.828 ;
      RECT 1.908 0.476 1.98 0.828 ;
      RECT 0.072 0.108 0.252 0.18 ;
      RECT 0.288 0.756 1.568 0.828 ;
      RECT 1.208 0.3 1.28 0.828 ;
      RECT 0.288 0.484 0.36 0.828 ;
      RECT 0.396 0.108 0.92 0.18 ;
  END
END XOR2x2_ASAP7_75t_R

MACRO XOR2xp5_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2xp5_ASAP7_75t_R 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.756 1.44 0.828 ;
        RECT 1.368 0.48 1.44 0.828 ;
        RECT 0.072 0.9 0.9 0.972 ;
        RECT 0.828 0.756 0.9 0.972 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.136 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.424 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.692 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.024 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.648 0.108 0.72 0.78 ;
      RECT 1.584 0.252 1.656 0.596 ;
      RECT 0.648 0.252 1.656 0.324 ;
      RECT 0.376 0.108 0.72 0.18 ;
      RECT 1.024 0.9 1.548 0.972 ;
  END
END XOR2xp5_ASAP7_75t_R

END LIBRARY ;

