../../libs/asap_7nm/asap7sc7p5t.datc_rdf.lef