asap7sc7p5t.datc_rdf.lef